module FFT8(clk, rst, i0, i1, i2, i3, i4, i5, i6, i7,
                o0, o1, o2, o3, o4, o5, o6, o7);
input clk, rst;
input [63:0] i0, i1, i2, i3, i4, i5, i6, i7;
output [63:0] o0, o1, o2, o3, o4, o5, o6, o7;
//---------------------------------------------------------------------------------
reg [63:0] o0, o1, o2, o3, o4, o5, o6, o7;

reg [31:0] sub1_0, sub1_1, sub1_2, sub1_3,
           sub2_0, sub2_1, sub2_2, sub2_3,
           sub2_c0, sub2_c1, sub2_c2, sub2_c3;
reg [64:0] real_0, real_1, real_2, real_3,
           imag_0, imag_1, imag_2, imag_3;
//---------------------------------------------------------------------------------
always@(posedge clk or posedge rst) begin
    if(rst) begin
        o0 = 0; o1 = 0; o2 = 0; o3 = 0;
        o4 = 0; o5 = 0; o6 = 0; o7 = 0;
    end else begin
        o0 = {i0[63:32] + i4[63:32], i0[31:0] + i4[31:0]};
        o1 = {i1[63:32] + i5[63:32], i1[31:0] + i5[31:0]};
        o2 = {i2[63:32] + i6[63:32], i2[31:0] + i6[31:0]};
        o3 = {i3[63:32] + i7[63:32], i3[31:0] + i7[31:0]};

        sub1_0 = i0[63:32] - i4[63:32];
        sub2_0 = i0[31:0] - i4[31:0];
        sub2_c0 = 0 - sub2_0;
        real_0 = {{32{sub1_0[31]}}, sub1_0} * {32'h0000, 32'h00010000} + {{32{sub2_c0[31]}}, sub2_c0} * {32'h0000, 32'h00000000};
        imag_0 = {{32{sub1_0[31]}}, sub1_0} * {32'h0000, 32'h00000000} + {{32{sub2_0[31]}}, sub2_0} * {32'h0000, 32'h00010000};
        o4 = {real_0[47:16], imag_0[47:16]};

        sub1_1 = i1[63:32] - i5[63:32];
        sub2_1 = i1[31:0] - i5[31:0];
        sub2_c1 = 0 - sub2_1;
        real_1 = {{32{sub1_1[31]}}, sub1_1} * {32'h0000, 32'h0000B504} + {{32{sub2_c1[31]}}, sub2_c1} * {32'hFFFF, 32'hFFFF4AFC};
        imag_1 = {{32{sub1_1[31]}}, sub1_1} * {32'hFFFF, 32'hFFFF4AFC} + {{32{sub2_1[31]}}, sub2_1} * {32'h0000, 32'h0000B504};
        o5 = {real_1[47:16], imag_1[47:16]};

        sub1_2 = i2[63:32] - i6[63:32];
        sub2_2 = i2[31:0] - i6[31:0];
        sub2_c2 = 0 - sub2_2;
        real_2 = {{32{sub1_2[31]}}, sub1_2} * {32'h0000, 32'h00000000} + {{32{sub2_c2[31]}}, sub2_c2} * {32'hFFFF, 32'hFFFF0000};
        imag_2 = {{32{sub1_2[31]}}, sub1_2} * {32'hFFFF, 32'hFFFF0000} + {{32{sub2_2[31]}}, sub2_2} * {32'h0000, 32'h00000000};
        o6 = {real_2[47:16], imag_2[47:16]};

        sub1_3 = i3[63:32] - i7[63:32];
        sub2_3 = i3[31:0] - i7[31:0];
        sub2_c3 = 0 - sub2_3;
        real_3 = {{32{sub1_3[31]}}, sub1_3} * {32'hFFFF, 32'hFFFF4AFC} + {{32{sub2_c3[31]}}, sub2_c3} * {32'hFFFF, 32'hFFFF4AFC};
        imag_3 = {{32{sub1_3[31]}}, sub1_3} * {32'hFFFF, 32'hFFFF4AFC} + {{32{sub2_3[31]}}, sub2_3} * {32'hFFFF, 32'hFFFF4AFC};
        o7 = {real_3[47:16], imag_3[47:16]};
    end
end

//---------------------------------------------------------------------------------
endmodule