module FFT16(clk, rst, i0, i1, i2, i3, i4, i5, i6, i7,
             i8, i9, ,i10 , i11, i12, i13, i14, i15,
             o0, o1, o2, o3, o4, o5, o6, o7, o8,
             o9, ,o10 , o11, o12, o13, o14, o15);
input clk, rst;
input [15:0] i0, i1, i2, i3, i4, i5, i6, i7, i8,
             i9, i10 , i11, i12, i13, i14, i15;
output [63:0] o0, o1, o2, o3, o4, o5, o6, o7, o8,
              o9, o10 , o11, o12, o13, o14, o15;
//---------------------------------------------------------------------------------
reg [63:0] o0, o1, o2, o3, o4, o5, o6, o7, o8,
            o9, o10 , o11, o12, o13, o14, o15;

reg [31:0] sub0, sub1, sub2, sub3, sub4, sub5, sub6, sub7;
reg [63:0] real_0, real_1, real_2, real_3, real_4, real_5, real_6, real_7,
           imag_0, imag_1, imag_2, imag_3, imag_4, imag_5, imag_6, imag_7;
//---------------------------------------------------------------------------------
always@(posedge clk or posedge rst) begin
    if(rst) begin
        o0 = 0; o1 = 0; o2 = 0; o3 = 0;
        o4 = 0; o5 = 0; o6 = 0; o7 = 0;
        o8 = 0; o9 = 0; o10 = 0; o11 = 0;
        o12 = 0; o13 = 0; o14 = 0; o15 = 0;
    end else begin
        o0 = {{{8{i0[15]}}, i0, 8'h00} + {{8{i8[15]}}, i8, 8'h00}, 32'h0000};
        o1 = {{{8{i1[15]}}, i1, 8'h00} + {{8{i9[15]}}, i9, 8'h00}, 32'h0000};
        o2 = {{{8{i2[15]}}, i2, 8'h00} + {{8{i10[15]}}, i10, 8'h00}, 32'h0000};
        o3 = {{{8{i3[15]}}, i3, 8'h00} + {{8{i11[15]}}, i11, 8'h00}, 32'h0000};
        o4 = {{{8{i4[15]}}, i4, 8'h00} + {{8{i12[15]}}, i12, 8'h00}, 32'h0000};
        o5 = {{{8{i5[15]}}, i5, 8'h00} + {{8{i13[15]}}, i13, 8'h00}, 32'h0000};
        o6 = {{{8{i6[15]}}, i6, 8'h00} + {{8{i14[15]}}, i14, 8'h00}, 32'h0000};
        o7 = {{{8{i7[15]}}, i7, 8'h00} + {{8{i15[15]}}, i15, 8'h00}, 32'h0000};

        sub0 = {{8{i0[15]}}, i0, 8'h00} - {{8{i8[15]}}, i8, 8'h00};
        real_0 = {{32{sub0[31]}}, sub0} * {32'h0000, 32'h00010000};
        imag_0 = {{32{sub0[31]}}, sub0} * {32'h0000, 32'h00000000};
        o8 = {real_0[47:16], imag_0[47:16]};

        sub1 = {{8{i1[15]}}, i1, 8'h00} - {{8{i9[15]}}, i9, 8'h00};
        real_1 = {{32{sub1[31]}}, sub1} * {32'h0000, 32'h0000EC83};
        imag_1 = {{32{sub1[31]}}, sub1} * {32'hFFFF, 32'hFFFF9E09};
        o9 = {real_1[47:16], imag_1[47:16]};

        sub2 = {{8{i2[15]}}, i2, 8'h00} - {{8{i10[15]}}, i10, 8'h00};
        real_2 = {{32{sub2[31]}}, sub2} * {32'h0000, 32'h0000B504};
        imag_2 = {{32{sub2[31]}}, sub2} * {32'hFFFF, 32'hFFFF4AFC};
        o10 = {real_2[47:16], imag_2[47:16]};

        sub3 = {{8{i3[15]}}, i3, 8'h00} - {{8{i11[15]}}, i11, 8'h00};
        real_3 = {{32{sub3[31]}}, sub3} * {32'h0000, 32'h000061F7};
        imag_3 = {{32{sub3[31]}}, sub3} * {32'hFFFF, 32'hFFFF137D};
        o11 = {real_3[47:16], imag_3[47:16]};

        sub4 = {{8{i4[15]}}, i4, 8'h00} - {{8{i12[15]}}, i12, 8'h00};
        real_4 = {{32{sub4[31]}}, sub4} * {32'h0000, 32'h00000000};
        imag_4 = {{32{sub4[31]}}, sub4} * {32'hFFFF, 32'hFFFF0000};
        o12 = {real_4[47:16], imag_4[47:16]};

        sub5 = {{8{i5[15]}}, i5, 8'h00} - {{8{i13[15]}}, i13, 8'h00};
        real_5 = {{32{sub5[31]}}, sub5} * {32'hFFFF, 32'hFFFF9E09};
        imag_5 = {{32{sub5[31]}}, sub5} * {32'hFFFF, 32'hFFFF137D};
        o13 = {real_5[47:16], imag_5[47:16]};

        sub6 = {{8{i6[15]}}, i6, 8'h00} - {{8{i14[15]}}, i14, 8'h00};
        real_6 = {{32{sub6[31]}}, sub6} * {32'hFFFF, 32'hFFFF4AFC};
        imag_6 = {{32{sub6[31]}}, sub6} * {32'hFFFF, 32'hFFFF4AFC};
        o14 = {real_6[47:16], imag_6[47:16]};

        sub7 = {{8{i7[15]}}, i7, 8'h00} - {{8{i15[15]}}, i15, 8'h00};
        real_7 = {{32{sub7[31]}}, sub7} * {32'hFFFF, 32'hFFFF137D};
        imag_7 = {{32{sub7[31]}}, sub7} * {32'hFFFF, 32'hFFFF9E09};
        o15 = {real_7[47:16], imag_7[47:16]};
    end
end

//---------------------------------------------------------------------------------
endmodule